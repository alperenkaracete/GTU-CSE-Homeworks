module slt_32bit(

input [31:0]A,
input [31:0]B,
output [31:0]Result
);

wire [31:0]notA;
wire [31:0]notB;
wire [31:0]or1;
wire [31:0]or2;

not notA1(notA[0],A[0]),
    notA2(notA[1],A[1]),
    notA3(notA[2],A[2]),
    notA4(notA[3],A[3]),
    notA5(notA[4],A[4]),
    notA6(notA[5],A[5]),
    notA7(notA[6],A[6]),
    notA8(notA[7],A[7]),
    notA9(notA[8],A[8]),
    notA10(notA[9],A[9]),
    notA11(notA[10],A[10]),
    notA12(notA[11],A[11]),
    notA13(notA[12],A[12]),
    notA14(notA[13],A[13]),
    notA15(notA[14],A[14]),
    notA16(notA[15],A[15]),
    notA17(notA[16],A[16]),
    notA18(notA[17],A[17]),
    notA19(notA[18],A[18]),
    notA20(notA[19],A[19]),
    notA21(notA[20],A[20]),
    notA22(notA[21],A[21]),
    notA23(notA[22],A[22]),
    notA24(notA[23],A[23]),
    notA25(notA[24],A[24]),
    notA26(notA[25],A[25]),
    notA27(notA[26],A[26]),
    notA28(notA[27],A[27]),
    notA29(notA[28],A[28]),
    notA30(notA[29],A[29]),
    notA31(notA[30],A[30]),
    notA32(notA[31],A[31]);

not notB1(notB[0],B[0]),
    notB2(notB[1],B[1]),
    notB3(notB[2],B[2]),
    notB4(notB[3],B[3]),
    notB5(notB[4],B[4]),
    notB6(notB[5],B[5]),
    notB7(notB[6],B[6]),
    notB8(notB[7],B[7]),
    notB9(notB[8],B[8]),
    notB10(notB[9],B[9]),
    notB11(notB[10],B[10]),
    notB12(notB[11],B[11]),
    notB13(notB[12],B[12]),
    notB14(notB[13],B[13]),
    notB15(notB[14],B[14]),
    notB16(notB[15],B[15]),
    notB17(notB[16],B[16]),
    notB18(notB[17],B[17]),
    notB19(notB[18],B[18]),
    notB20(notB[19],B[19]),
    notB21(notB[20],B[20]),
    notB22(notB[21],B[21]),
    notB23(notB[22],B[22]),
    notB24(notB[23],B[23]),
    notB25(notB[24],B[24]),
    notB26(notB[25],B[25]),
    notB27(notB[26],B[26]),
    notB28(notB[27],B[27]),
    notB29(notB[28],B[28]),
    notB30(notB[29],B[29]),
    notB31(notB[30],B[30]),
    notB32(notB[31],B[31]);  
    
or  orA1(or1[0],notA[0],B[0]),
    orA2(or1[1],notA[1],B[1]),
    orA3(or1[2],notA[2],B[2]),
    orA4(or1[3],notA[3],B[3]),
    orA5(or1[4],notA[4],B[4]),
    orA6(or1[5],notA[5],B[5]),
    orA7(or1[6],notA[6],B[6]),
    orA8(or1[7],notA[7],B[7]),
    orA9(or1[8],notA[8],B[8]),
    orA10(or1[9],notA[9],B[9]),
    orA11(or1[10],notA[10],B[10]),
    orA12(or1[11],notA[11],B[11]),
    orA13(or1[12],notA[12],B[12]),
    orA14(or1[13],notA[13],B[13]),
    orA15(or1[14],notA[14],B[14]),
    orA16(or1[15],notA[15],B[15]),
    orA17(or1[16],notA[16],B[16]),
    orA18(or1[17],notA[17],B[17]),
    orA19(or1[18],notA[18],B[18]),
    orA20(or1[19],notA[19],B[19]),
    orA21(or1[20],notA[20],B[20]),
    orA22(or1[21],notA[21],B[21]),
    orA23(or1[22],notA[22],B[22]),
    orA24(or1[23],notA[23],B[23]),
    orA25(or1[24],notA[24],B[24]),
    orA26(or1[25],notA[25],B[25]),
    orA27(or1[26],notA[26],B[26]),
    orA28(or1[27],notA[27],B[27]),
    orA29(or1[28],notA[28],B[28]),
    orA30(or1[29],notA[29],B[29]),
    orA31(or1[30],notA[30],B[30]),
    orA32(or1[31],notA[31],B[31]); 

or  orB1(or2[0],notB[0],A[0]),
    orB2(or2[1],notB[1],A[1]),
    orB3(or2[2],notB[2],A[2]),
    orB4(or2[3],notB[3],A[3]),
    orB5(or2[4],notB[4],A[4]),
    orB6(or2[5],notB[5],A[5]),
    orB7(or2[6],notB[6],A[6]),
    orB8(or2[7],notB[7],A[7]),
    orB9(or2[8],notB[8],A[8]),
    orB10(or2[9],notB[9],A[9]),
    orB11(or2[10],notB[10],A[10]),
    orB12(or2[11],notB[11],A[11]),
    orB13(or2[12],notB[12],A[12]),
    orB14(or2[13],notB[13],A[13]),
    orB15(or2[14],notB[14],A[14]),
    orB16(or2[15],notB[15],A[15]),
    orB17(or2[16],notB[16],A[16]),
    orB18(or2[17],notB[17],A[17]),
    orB19(or2[18],notB[18],A[18]),
    orB20(or2[19],notB[19],A[19]),
    orB21(or2[20],notB[20],A[20]),
    orB22(or2[21],notB[21],A[21]),
    orB23(or2[22],notB[22],A[22]),
    orB24(or2[23],notB[23],A[23]),
    orB25(or2[24],notB[24],A[24]),
    orB26(or2[25],notB[25],A[25]),
    orB27(or2[26],notB[26],A[26]),
    orB28(or2[27],notB[27],A[27]),
    orB29(or2[28],notB[28],A[28]),
    orB30(or2[29],notB[29],A[29]),
    orB31(or2[30],notB[30],A[30]),
    orB32(or2[31],notB[31],A[31]);     

and and1(Result[0],or1[0],or2[0]),
    and2(Result[1],or1[1],or2[1]),
    and3(Result[2],or1[2],or2[2]),
    and4(Result[3],or1[3],or2[3]),
    and5(Result[4],or1[4],or2[4]),
    and6(Result[5],or1[5],or2[5]),
    and7(Result[6],or1[6],or2[6]),
    and8(Result[7],or1[7],or2[7]),
    and9(Result[8],or1[8],or2[8]),
    and10(Result[9],or1[9],or2[9]),
    and11(Result[10],or1[10],or2[10]),
    and12(Result[11],or1[11],or2[11]),
    and13(Result[12],or1[12],or2[12]),
    and14(Result[13],or1[13],or2[13]),
    and15(Result[14],or1[14],or2[14]),
    and16(Result[15],or1[15],or2[15]),
    and17(Result[16],or1[16],or2[16]),
    and18(Result[17],or1[17],or2[17]),
    and19(Result[18],or1[18],or2[18]),
    and20(Result[19],or1[19],or2[19]),
    and21(Result[20],or1[20],or2[20]),
    and22(Result[21],or1[21],or2[21]),
    and23(Result[22],or1[22],or2[22]),
    and24(Result[23],or1[23],or2[23]),
    and25(Result[24],or1[24],or2[24]),
    and26(Result[25],or1[25],or2[25]),
    and27(Result[26],or1[26],or2[26]),
    and28(Result[27],or1[27],or2[27]),
    and29(Result[28],or1[28],or2[28]),
    and30(Result[29],or1[29],or2[29]),
    and31(Result[30],or1[30],or2[30]),
    and32(Result[31],or1[31],or2[31]);
	 
endmodule
